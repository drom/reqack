// edge ${id} EB1
always @(posedge clk) if (en_${id}) ${i_0_data} <= ${t_0_data};
